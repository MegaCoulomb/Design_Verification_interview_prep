// TODO: Build UVM testbench for arbiter
