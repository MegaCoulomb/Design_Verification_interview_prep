// TODO: Build UVM testbench for cache
