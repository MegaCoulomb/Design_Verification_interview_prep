class fifo_scoreboard extends uvm_component;
  `uvm_component_utils(fifo_scoreboard)
  function new(string name, uvm_component parent); super.new(name,parent); endfunction
endclass
