// TODO: Implement 3‑stage pipelined CPU
