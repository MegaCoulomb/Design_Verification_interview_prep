// TODO: FPGA top‑level integration wrapper
