// TODO: CPU verification env
