// TODO: Implement fair round‑robin arbiter
