// TODO: Implement direct‑mapped cache
