`ifndef UVM_INCLUDES_SVH
`define UVM_INCLUDES_SVH
`include "uvm_macros.svh"
import uvm_pkg::*;
`endif
